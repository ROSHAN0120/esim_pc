* D:\eSim_tut\files\PC\PC.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 05/26/23 22:26:18

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U10  1 2 3 4 5 6 7 8 Net-_U10-Pad9_ Net-_U10-Pad10_ Net-_U10-Pad11_ Net-_U10-Pad12_ Net-_U10-Pad13_ Net-_U10-Pad14_ Net-_U10-Pad15_ Net-_U10-Pad16_ adc_bridge_8		
U11  Net-_U11-Pad1_ Net-_U11-Pad2_ Net-_U11-Pad3_ Net-_U11-Pad4_ o1 o2 o3 o4 dac_bridge_4		
v1  1 GND pulse		
v2  2 GND pulse		
v3  3 GND pulse		
v4  4 GND pulse		
v5  5 GND pulse		
v6  6 GND pulse		
v7  7 GND pulse		
v8  8 GND pulse		
U6  3 plot_v1		
U8  4 plot_v1		
U9  5 plot_v1		
U7  6 plot_v1		
U5  7 plot_v1		
U2  8 plot_v1		
U1  1 plot_v1		
U4  2 plot_v1		
U13  o3 plot_v1		
U12  o4 plot_v1		
U15  o1 plot_v1		
U14  o2 plot_v1		
U3  Net-_U10-Pad9_ Net-_U10-Pad10_ Net-_U10-Pad11_ Net-_U10-Pad12_ Net-_U10-Pad13_ Net-_U10-Pad14_ Net-_U10-Pad15_ Net-_U10-Pad16_ Net-_U11-Pad1_ Net-_U11-Pad2_ Net-_U11-Pad3_ Net-_U11-Pad4_ pc		

.end
